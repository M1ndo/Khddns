module main

import args

fn main() {
	args.parser()!
}
